module desloca2(input logic [31:0] a, output logic [31:0] s);

assign s = a << 2;

endmodule